`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/05/09 20:36:21
// Design Name: 
// Module Name: MULT
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MULT(
    input [31:0] a,
    input [31:0] b,
    output [31:0] hi,
    output [31:0] lo
    );
    wire [63:0] moved_a[31:0];
    wire [63:0] z;
    assign moved_a[0]=(b[0])?(-{{32{a[31]}},a}):64'b0;
    assign moved_a[1]=(b[1]^b[0])?(b[1]?(-{{31{a[31]}},a,1'b0}):({{31{a[31]}},a,1'b0})):64'b0;
    assign moved_a[2]=(b[2]^b[1])?(b[2]?(-{{30{a[31]}},a,2'b0}):({{30{a[31]}},a,2'b0})):64'b0;
    assign moved_a[3]=(b[3]^b[2])?(b[3]?(-{{29{a[31]}},a,3'b0}):({{29{a[31]}},a,3'b0})):64'b0;
    assign moved_a[4]=(b[4]^b[3])?(b[4]?(-{{28{a[31]}},a,4'b0}):({{28{a[31]}},a,4'b0})):64'b0;
    assign moved_a[5]=(b[5]^b[4])?(b[5]?(-{{27{a[31]}},a,5'b0}):({{27{a[31]}},a,5'b0})):64'b0;
    assign moved_a[6]=(b[6]^b[5])?(b[6]?(-{{26{a[31]}},a,6'b0}):({{26{a[31]}},a,6'b0})):64'b0;
    assign moved_a[7]=(b[7]^b[6])?(b[7]?(-{{25{a[31]}},a,7'b0}):({{25{a[31]}},a,7'b0})):64'b0;
    assign moved_a[8]=(b[8]^b[7])?(b[8]?(-{{24{a[31]}},a,8'b0}):({{24{a[31]}},a,8'b0})):64'b0;
    assign moved_a[9]=(b[9]^b[8])?(b[9]?(-{{23{a[31]}},a,9'b0}):({{23{a[31]}},a,9'b0})):64'b0;
    assign moved_a[10]=(b[10]^b[9])?(b[10]?(-{{22{a[31]}},a,10'b0}):({{22{a[31]}},a,10'b0})):64'b0;
    assign moved_a[11]=(b[11]^b[10])?(b[11]?(-{{21{a[31]}},a,11'b0}):({{21{a[31]}},a,11'b0})):64'b0;
    assign moved_a[12]=(b[12]^b[11])?(b[12]?(-{{20{a[31]}},a,12'b0}):({{20{a[31]}},a,12'b0})):64'b0;
    assign moved_a[13]=(b[13]^b[12])?(b[13]?(-{{19{a[31]}},a,13'b0}):({{19{a[31]}},a,13'b0})):64'b0;
    assign moved_a[14]=(b[14]^b[13])?(b[14]?(-{{18{a[31]}},a,14'b0}):({{18{a[31]}},a,14'b0})):64'b0;
    assign moved_a[15]=(b[15]^b[14])?(b[15]?(-{{17{a[31]}},a,15'b0}):({{17{a[31]}},a,15'b0})):64'b0;
    assign moved_a[16]=(b[16]^b[15])?(b[16]?(-{{16{a[31]}},a,16'b0}):({{16{a[31]}},a,16'b0})):64'b0;
    assign moved_a[17]=(b[17]^b[16])?(b[17]?(-{{15{a[31]}},a,17'b0}):({{15{a[31]}},a,17'b0})):64'b0;
    assign moved_a[18]=(b[18]^b[17])?(b[18]?(-{{14{a[31]}},a,18'b0}):({{14{a[31]}},a,18'b0})):64'b0;
    assign moved_a[19]=(b[19]^b[18])?(b[19]?(-{{13{a[31]}},a,19'b0}):({{13{a[31]}},a,19'b0})):64'b0;
    assign moved_a[20]=(b[20]^b[19])?(b[20]?(-{{12{a[31]}},a,20'b0}):({{12{a[31]}},a,20'b0})):64'b0;
    assign moved_a[21]=(b[21]^b[20])?(b[21]?(-{{11{a[31]}},a,21'b0}):({{11{a[31]}},a,21'b0})):64'b0;
    assign moved_a[22]=(b[22]^b[21])?(b[22]?(-{{10{a[31]}},a,22'b0}):({{10{a[31]}},a,22'b0})):64'b0;
    assign moved_a[23]=(b[23]^b[22])?(b[23]?(-{{9{a[31]}},a,23'b0}):({{9{a[31]}},a,23'b0})):64'b0;
    assign moved_a[24]=(b[24]^b[23])?(b[24]?(-{{8{a[31]}},a,24'b0}):({{8{a[31]}},a,24'b0})):64'b0;
    assign moved_a[25]=(b[25]^b[24])?(b[25]?(-{{7{a[31]}},a,25'b0}):({{7{a[31]}},a,25'b0})):64'b0;
    assign moved_a[26]=(b[26]^b[25])?(b[26]?(-{{6{a[31]}},a,26'b0}):({{6{a[31]}},a,26'b0})):64'b0;
    assign moved_a[27]=(b[27]^b[26])?(b[27]?(-{{5{a[31]}},a,27'b0}):({{5{a[31]}},a,27'b0})):64'b0;
    assign moved_a[28]=(b[28]^b[27])?(b[28]?(-{{4{a[31]}},a,28'b0}):({{4{a[31]}},a,28'b0})):64'b0;
    assign moved_a[29]=(b[29]^b[28])?(b[29]?(-{{3{a[31]}},a,29'b0}):({{3{a[31]}},a,29'b0})):64'b0;
    assign moved_a[30]=(b[30]^b[29])?(b[30]?(-{{2{a[31]}},a,30'b0}):({{2{a[31]}},a,30'b0})):64'b0;
    assign moved_a[31]=(b[31]^b[30])?(b[31]?(-{{1{a[31]}},a,31'b0}):({{1{a[31]}},a,31'b0})):64'b0;
    assign z=moved_a[0]+moved_a[1]+moved_a[2]+moved_a[3]+moved_a[4]
            +moved_a[5]+moved_a[6]+moved_a[7]+moved_a[8]+moved_a[9]
            +moved_a[10]+moved_a[11]+moved_a[12]+moved_a[13]+moved_a[14]
            +moved_a[15]+moved_a[16]+moved_a[17]+moved_a[18]+moved_a[19]
            +moved_a[20]+moved_a[21]+moved_a[22]+moved_a[23]+moved_a[24]
            +moved_a[25]+moved_a[26]+moved_a[27]+moved_a[28]+moved_a[29]
            +moved_a[30]+moved_a[31];
    assign hi=z[63:32];
    assign lo=z[31:0];
endmodule
